magic
tech scmos
timestamp 1731952171
<< nwell >>
rect 371 367 429 391
rect 444 335 511 391
rect 527 367 552 391
rect 558 335 604 391
rect 621 367 679 391
rect 383 267 407 294
rect 422 237 446 264
rect 556 245 599 269
rect 633 267 657 294
rect 672 237 696 264
rect 386 184 488 208
rect 520 184 545 208
rect 551 168 583 208
rect 595 184 653 208
rect 434 110 450 134
rect 459 115 486 139
rect 397 83 421 110
rect 537 75 580 99
rect 607 84 631 111
rect 646 54 670 81
<< ntransistor >>
rect 384 356 386 359
rect 415 356 417 359
rect 538 356 540 359
rect 634 356 636 359
rect 665 356 667 359
rect 368 328 374 330
rect 383 328 389 330
rect 408 328 414 330
rect 423 328 429 330
rect 618 328 624 330
rect 633 328 639 330
rect 658 328 664 330
rect 673 328 679 330
rect 368 306 374 308
rect 383 306 389 308
rect 526 320 532 322
rect 541 320 547 322
rect 485 315 487 318
rect 583 316 585 319
rect 408 306 414 308
rect 423 306 429 308
rect 477 307 479 310
rect 493 307 495 310
rect 575 308 577 311
rect 591 308 593 311
rect 618 306 624 308
rect 633 306 639 308
rect 658 306 664 308
rect 673 306 679 308
rect 469 292 471 295
rect 485 292 487 295
rect 501 292 503 295
rect 567 293 569 296
rect 583 293 585 296
rect 599 293 601 296
rect 372 279 375 281
rect 622 279 625 281
rect 477 269 479 272
rect 493 269 495 272
rect 411 249 414 251
rect 661 249 664 251
rect 569 234 571 237
rect 585 234 587 237
rect 399 173 401 176
rect 430 173 432 176
rect 458 173 460 176
rect 474 173 476 176
rect 531 173 533 176
rect 608 173 610 176
rect 639 173 641 176
rect 383 145 389 147
rect 398 145 404 147
rect 423 145 429 147
rect 438 145 444 147
rect 565 148 567 151
rect 592 145 598 147
rect 607 145 613 147
rect 632 145 638 147
rect 647 145 653 147
rect 557 140 559 143
rect 573 140 575 143
rect 519 137 525 139
rect 534 137 540 139
rect 423 121 426 123
rect 592 123 598 125
rect 607 123 613 125
rect 632 123 638 125
rect 647 123 653 125
rect 497 108 499 114
rect 472 104 474 107
rect 386 95 389 97
rect 497 93 499 99
rect 596 96 599 98
rect 550 64 552 67
rect 566 64 568 67
rect 635 66 638 68
<< ptransistor >>
rect 384 373 386 384
rect 415 373 417 384
rect 480 378 484 380
rect 538 373 540 384
rect 564 378 568 380
rect 466 370 470 372
rect 496 370 500 372
rect 452 362 456 364
rect 476 362 480 364
rect 634 373 636 384
rect 665 373 667 384
rect 578 370 582 372
rect 568 362 572 364
rect 592 362 596 364
rect 466 354 470 356
rect 496 354 500 356
rect 578 354 582 356
rect 480 346 484 348
rect 568 346 572 348
rect 389 279 400 281
rect 639 279 650 281
rect 428 249 439 251
rect 569 251 571 262
rect 585 251 587 262
rect 678 249 689 251
rect 399 190 401 201
rect 430 190 432 201
rect 458 190 460 201
rect 474 190 476 201
rect 531 190 533 201
rect 561 195 565 197
rect 608 190 610 201
rect 639 190 641 201
rect 571 187 575 189
rect 557 179 561 181
rect 440 121 444 123
rect 472 121 474 132
rect 403 95 414 97
rect 613 96 624 98
rect 550 81 552 92
rect 566 81 568 92
rect 652 66 663 68
<< ndiffusion >>
rect 383 356 384 359
rect 386 356 387 359
rect 414 356 415 359
rect 417 356 418 359
rect 537 356 538 359
rect 540 356 541 359
rect 633 356 634 359
rect 636 356 637 359
rect 664 356 665 359
rect 667 356 668 359
rect 368 330 374 331
rect 383 330 389 331
rect 408 330 414 331
rect 423 330 429 331
rect 618 330 624 331
rect 633 330 639 331
rect 658 330 664 331
rect 673 330 679 331
rect 368 327 374 328
rect 383 327 389 328
rect 408 327 414 328
rect 423 327 429 328
rect 618 327 624 328
rect 368 308 374 309
rect 383 308 389 309
rect 408 308 414 309
rect 423 308 429 309
rect 526 322 532 323
rect 541 322 547 323
rect 484 315 485 318
rect 487 315 488 318
rect 526 319 532 320
rect 541 319 547 320
rect 633 327 639 328
rect 658 327 664 328
rect 673 327 679 328
rect 582 316 583 319
rect 585 316 586 319
rect 476 307 477 310
rect 479 307 480 310
rect 492 307 493 310
rect 495 307 496 310
rect 574 308 575 311
rect 577 308 578 311
rect 590 308 591 311
rect 593 308 594 311
rect 618 308 624 309
rect 633 308 639 309
rect 368 305 374 306
rect 383 305 389 306
rect 408 305 414 306
rect 423 305 429 306
rect 658 308 664 309
rect 673 308 679 309
rect 618 305 624 306
rect 633 305 639 306
rect 658 305 664 306
rect 673 305 679 306
rect 468 292 469 295
rect 471 292 472 295
rect 372 281 375 282
rect 484 292 485 295
rect 487 292 488 295
rect 500 292 501 295
rect 503 292 504 295
rect 566 293 567 296
rect 569 293 570 296
rect 582 293 583 296
rect 585 293 586 296
rect 598 293 599 296
rect 601 293 602 296
rect 372 278 375 279
rect 622 281 625 282
rect 622 278 625 279
rect 476 269 477 272
rect 479 269 480 272
rect 492 269 493 272
rect 495 269 496 272
rect 411 251 414 252
rect 411 248 414 249
rect 661 251 664 252
rect 661 248 664 249
rect 568 234 569 237
rect 571 234 572 237
rect 584 234 585 237
rect 587 234 588 237
rect 398 173 399 176
rect 401 173 402 176
rect 429 173 430 176
rect 432 173 433 176
rect 457 173 458 176
rect 460 173 461 176
rect 473 173 474 176
rect 476 173 477 176
rect 530 173 531 176
rect 533 173 534 176
rect 607 173 608 176
rect 610 173 611 176
rect 638 173 639 176
rect 641 173 642 176
rect 383 147 389 148
rect 398 147 404 148
rect 423 147 429 148
rect 438 147 444 148
rect 383 144 389 145
rect 398 144 404 145
rect 423 144 429 145
rect 438 144 444 145
rect 564 148 565 151
rect 567 148 568 151
rect 592 147 598 148
rect 607 147 613 148
rect 632 147 638 148
rect 647 147 653 148
rect 592 144 598 145
rect 519 139 525 140
rect 556 140 557 143
rect 559 140 560 143
rect 572 140 573 143
rect 575 140 576 143
rect 607 144 613 145
rect 632 144 638 145
rect 647 144 653 145
rect 534 139 540 140
rect 519 136 525 137
rect 534 136 540 137
rect 423 123 426 124
rect 423 120 426 121
rect 592 125 598 126
rect 607 125 613 126
rect 632 125 638 126
rect 647 125 653 126
rect 592 122 598 123
rect 607 122 613 123
rect 632 122 638 123
rect 647 122 653 123
rect 496 108 497 114
rect 499 108 500 114
rect 471 104 472 107
rect 474 104 475 107
rect 386 97 389 98
rect 386 94 389 95
rect 496 93 497 99
rect 499 93 500 99
rect 596 98 599 99
rect 596 95 599 96
rect 635 68 638 69
rect 549 64 550 67
rect 552 64 553 67
rect 565 64 566 67
rect 568 64 569 67
rect 635 65 638 66
<< pdiffusion >>
rect 383 373 384 384
rect 386 373 387 384
rect 414 373 415 384
rect 417 373 418 384
rect 480 380 484 381
rect 480 377 484 378
rect 466 372 470 373
rect 496 372 500 373
rect 537 373 538 384
rect 540 373 541 384
rect 564 380 568 381
rect 564 377 568 378
rect 466 369 470 370
rect 496 369 500 370
rect 452 364 456 365
rect 476 364 480 365
rect 452 361 456 362
rect 476 361 480 362
rect 466 356 470 357
rect 496 356 500 357
rect 578 372 582 373
rect 633 373 634 384
rect 636 373 637 384
rect 664 373 665 384
rect 667 373 668 384
rect 578 369 582 370
rect 568 364 572 365
rect 592 364 596 365
rect 568 361 572 362
rect 592 361 596 362
rect 578 356 582 357
rect 466 353 470 354
rect 496 353 500 354
rect 578 353 582 354
rect 480 348 484 349
rect 568 348 572 349
rect 480 345 484 346
rect 568 345 572 346
rect 389 281 400 282
rect 389 278 400 279
rect 639 281 650 282
rect 639 278 650 279
rect 428 251 439 252
rect 428 248 439 249
rect 568 251 569 262
rect 571 251 572 262
rect 584 251 585 262
rect 587 251 588 262
rect 678 251 689 252
rect 678 248 689 249
rect 398 190 399 201
rect 401 190 402 201
rect 429 190 430 201
rect 432 190 433 201
rect 457 190 458 201
rect 460 190 461 201
rect 473 190 474 201
rect 476 190 477 201
rect 530 190 531 201
rect 533 190 534 201
rect 561 197 565 198
rect 561 194 565 195
rect 607 190 608 201
rect 610 190 611 201
rect 638 190 639 201
rect 641 190 642 201
rect 571 189 575 190
rect 571 186 575 187
rect 557 181 561 182
rect 557 178 561 179
rect 440 123 444 124
rect 440 120 444 121
rect 471 121 472 132
rect 474 121 475 132
rect 403 97 414 98
rect 403 94 414 95
rect 613 98 624 99
rect 549 81 550 92
rect 552 81 553 92
rect 565 81 566 92
rect 568 81 569 92
rect 613 95 624 96
rect 652 68 663 69
rect 652 65 663 66
<< ndcontact >>
rect 379 355 383 359
rect 387 355 391 359
rect 410 355 414 359
rect 418 355 422 359
rect 533 355 537 359
rect 541 355 545 359
rect 629 355 633 359
rect 637 355 641 359
rect 660 355 664 359
rect 668 355 672 359
rect 368 331 374 335
rect 383 331 389 335
rect 408 331 414 335
rect 423 331 429 335
rect 618 331 624 335
rect 633 331 639 335
rect 658 331 664 335
rect 673 331 679 335
rect 368 323 374 327
rect 383 323 389 327
rect 408 323 414 327
rect 423 323 429 327
rect 368 309 374 313
rect 383 309 389 313
rect 408 309 414 313
rect 423 309 429 313
rect 480 315 484 319
rect 526 323 532 327
rect 541 323 547 327
rect 488 315 492 319
rect 526 315 532 319
rect 541 315 547 319
rect 578 316 582 320
rect 618 323 624 327
rect 633 323 639 327
rect 658 323 664 327
rect 673 323 679 327
rect 586 316 590 320
rect 472 307 476 311
rect 480 307 484 311
rect 488 307 492 311
rect 496 307 500 311
rect 570 308 574 312
rect 578 308 582 312
rect 586 308 590 312
rect 594 308 598 312
rect 618 309 624 313
rect 633 309 639 313
rect 368 301 374 305
rect 383 301 389 305
rect 408 301 414 305
rect 423 301 429 305
rect 658 309 664 313
rect 673 309 679 313
rect 618 301 624 305
rect 633 301 639 305
rect 658 301 664 305
rect 673 301 679 305
rect 464 291 468 295
rect 371 282 375 286
rect 472 291 476 295
rect 480 291 484 295
rect 488 291 492 295
rect 496 291 500 295
rect 504 291 508 295
rect 562 292 566 296
rect 570 292 574 296
rect 578 292 582 296
rect 586 292 590 296
rect 594 292 598 296
rect 602 292 606 296
rect 371 274 375 278
rect 621 282 625 286
rect 621 274 625 278
rect 472 268 476 272
rect 480 268 484 272
rect 488 268 492 272
rect 496 268 500 272
rect 410 252 414 256
rect 410 244 414 248
rect 660 252 664 256
rect 660 244 664 248
rect 564 233 568 237
rect 572 233 576 237
rect 580 233 584 237
rect 588 233 592 237
rect 394 172 398 176
rect 402 172 406 176
rect 425 172 429 176
rect 433 172 437 176
rect 453 172 457 176
rect 461 172 465 176
rect 469 172 473 176
rect 477 172 481 176
rect 526 172 530 176
rect 534 172 538 176
rect 603 172 607 176
rect 611 172 615 176
rect 634 172 638 176
rect 642 172 646 176
rect 383 148 389 152
rect 398 148 404 152
rect 423 148 429 152
rect 438 148 444 152
rect 383 140 389 144
rect 398 140 404 144
rect 423 140 429 144
rect 560 148 564 152
rect 568 148 572 152
rect 592 148 598 152
rect 607 148 613 152
rect 632 148 638 152
rect 647 148 653 152
rect 438 140 444 144
rect 519 140 525 144
rect 534 140 540 144
rect 552 140 556 144
rect 560 140 564 144
rect 568 140 572 144
rect 576 140 580 144
rect 592 140 598 144
rect 607 140 613 144
rect 632 140 638 144
rect 647 140 653 144
rect 519 132 525 136
rect 534 132 540 136
rect 422 124 426 128
rect 422 116 426 120
rect 592 126 598 130
rect 607 126 613 130
rect 632 126 638 130
rect 647 126 653 130
rect 592 118 598 122
rect 607 118 613 122
rect 632 118 638 122
rect 647 118 653 122
rect 492 108 496 114
rect 500 108 504 114
rect 467 103 471 107
rect 475 103 479 107
rect 385 98 389 102
rect 595 99 599 103
rect 385 90 389 94
rect 492 93 496 99
rect 500 93 504 99
rect 595 91 599 95
rect 634 69 638 73
rect 545 63 549 67
rect 553 63 557 67
rect 561 63 565 67
rect 569 63 573 67
rect 634 61 638 65
<< pdcontact >>
rect 379 373 383 384
rect 387 373 391 384
rect 410 373 414 384
rect 418 373 422 384
rect 480 381 484 385
rect 466 373 470 377
rect 480 373 484 377
rect 496 373 500 377
rect 533 373 537 384
rect 541 373 545 384
rect 564 381 568 385
rect 564 373 568 377
rect 578 373 582 377
rect 452 365 456 369
rect 466 365 470 369
rect 476 365 480 369
rect 496 365 500 369
rect 452 357 456 361
rect 466 357 470 361
rect 476 357 480 361
rect 496 357 500 361
rect 629 373 633 384
rect 637 373 641 384
rect 660 373 664 384
rect 668 373 672 384
rect 568 365 572 369
rect 578 365 582 369
rect 592 365 596 369
rect 568 357 572 361
rect 578 357 582 361
rect 592 357 596 361
rect 466 349 470 353
rect 480 349 484 353
rect 496 349 500 353
rect 568 349 572 353
rect 578 349 582 353
rect 480 341 484 345
rect 568 341 572 345
rect 389 282 400 286
rect 639 282 650 286
rect 389 274 400 278
rect 639 274 650 278
rect 428 252 439 256
rect 564 251 568 262
rect 572 251 576 262
rect 580 251 584 262
rect 588 251 592 262
rect 678 252 689 256
rect 428 244 439 248
rect 678 244 689 248
rect 394 190 398 201
rect 402 190 406 201
rect 425 190 429 201
rect 433 190 437 201
rect 453 190 457 201
rect 461 190 465 201
rect 469 190 473 201
rect 477 190 481 201
rect 526 190 530 201
rect 534 190 538 201
rect 561 198 565 202
rect 561 190 565 194
rect 571 190 575 194
rect 603 190 607 201
rect 611 190 615 201
rect 634 190 638 201
rect 642 190 646 201
rect 557 182 561 186
rect 571 182 575 186
rect 557 174 561 178
rect 440 124 444 128
rect 467 121 471 132
rect 475 121 479 132
rect 440 116 444 120
rect 403 98 414 102
rect 403 90 414 94
rect 613 99 624 103
rect 545 81 549 92
rect 553 81 557 92
rect 561 81 565 92
rect 569 81 573 92
rect 613 91 624 95
rect 652 69 663 73
rect 652 61 663 65
<< psubstratepcontact >>
rect 379 346 383 350
rect 410 346 414 350
rect 541 344 545 348
rect 629 346 633 350
rect 660 346 664 350
rect 361 281 365 285
rect 611 281 615 285
rect 399 252 403 256
rect 649 252 653 256
rect 564 222 568 226
rect 580 222 584 226
rect 394 162 398 166
rect 425 161 429 165
rect 461 161 465 165
rect 477 161 481 165
rect 534 161 538 165
rect 603 163 607 167
rect 634 163 638 167
rect 411 124 415 128
rect 564 131 568 135
rect 374 98 378 102
rect 584 99 588 103
rect 467 92 471 96
rect 623 69 627 73
rect 545 52 549 56
rect 561 52 565 56
<< nsubstratencontact >>
rect 383 391 387 395
rect 414 391 418 395
rect 472 391 476 395
rect 633 391 637 395
rect 664 391 668 395
rect 407 278 411 282
rect 657 278 661 282
rect 568 269 572 273
rect 584 269 588 273
rect 446 248 450 252
rect 696 248 700 252
rect 398 208 402 212
rect 429 208 433 212
rect 457 208 461 212
rect 473 208 477 212
rect 530 208 534 212
rect 564 208 568 212
rect 607 208 611 212
rect 638 208 642 212
rect 471 139 475 143
rect 450 120 454 124
rect 549 99 553 103
rect 565 99 569 103
rect 421 94 425 98
rect 631 95 635 99
rect 670 65 674 69
<< polysilicon >>
rect 384 384 386 387
rect 415 384 417 387
rect 538 384 540 387
rect 473 378 480 380
rect 484 378 487 380
rect 384 359 386 373
rect 415 359 417 373
rect 634 384 636 387
rect 665 384 667 387
rect 561 378 564 380
rect 568 378 575 380
rect 459 370 466 372
rect 470 370 473 372
rect 493 370 496 372
rect 500 370 507 372
rect 445 362 452 364
rect 456 362 459 364
rect 473 362 476 364
rect 480 362 487 364
rect 538 359 540 373
rect 575 370 578 372
rect 582 370 589 372
rect 561 362 568 364
rect 572 362 575 364
rect 589 362 592 364
rect 596 362 603 364
rect 384 351 386 355
rect 415 351 417 355
rect 459 354 466 356
rect 470 354 473 356
rect 493 354 496 356
rect 500 354 507 356
rect 634 359 636 373
rect 665 359 667 373
rect 538 351 540 355
rect 575 354 578 356
rect 582 354 589 356
rect 634 351 636 355
rect 665 351 667 355
rect 473 346 480 348
rect 484 346 487 348
rect 561 346 568 348
rect 572 346 575 348
rect 361 328 368 330
rect 374 328 377 330
rect 380 328 383 330
rect 389 328 396 330
rect 401 328 408 330
rect 414 328 417 330
rect 420 328 423 330
rect 429 328 436 330
rect 611 328 618 330
rect 624 328 627 330
rect 630 328 633 330
rect 639 328 646 330
rect 651 328 658 330
rect 664 328 667 330
rect 670 328 673 330
rect 679 328 686 330
rect 361 306 368 308
rect 374 306 377 308
rect 380 306 383 308
rect 389 306 396 308
rect 477 311 479 318
rect 485 318 487 326
rect 519 320 526 322
rect 532 320 535 322
rect 538 320 541 322
rect 547 320 554 322
rect 485 312 487 314
rect 493 311 495 318
rect 575 312 577 319
rect 583 319 585 327
rect 583 313 585 315
rect 591 312 593 319
rect 401 306 408 308
rect 414 306 417 308
rect 420 306 423 308
rect 429 306 436 308
rect 477 304 479 307
rect 493 304 495 307
rect 575 305 577 308
rect 591 305 593 308
rect 611 306 618 308
rect 624 306 627 308
rect 630 306 633 308
rect 639 306 646 308
rect 651 306 658 308
rect 664 306 667 308
rect 670 306 673 308
rect 679 306 686 308
rect 469 295 471 298
rect 485 295 487 298
rect 501 295 503 298
rect 567 296 569 299
rect 583 296 585 299
rect 599 296 601 299
rect 469 284 471 292
rect 485 284 487 292
rect 501 284 503 292
rect 567 285 569 293
rect 583 285 585 293
rect 599 285 601 293
rect 367 279 371 281
rect 375 279 389 281
rect 400 279 403 281
rect 617 279 621 281
rect 625 279 639 281
rect 650 279 653 281
rect 477 272 479 275
rect 493 272 495 275
rect 477 261 479 268
rect 493 261 495 268
rect 569 262 571 265
rect 585 262 587 265
rect 406 249 410 251
rect 414 249 428 251
rect 439 249 442 251
rect 569 237 571 251
rect 585 237 587 251
rect 656 249 660 251
rect 664 249 678 251
rect 689 249 692 251
rect 569 229 571 233
rect 585 229 587 233
rect 399 201 401 204
rect 430 201 432 204
rect 458 201 460 204
rect 474 201 476 204
rect 531 201 533 204
rect 608 201 610 204
rect 639 201 641 204
rect 554 195 561 197
rect 565 195 568 197
rect 399 176 401 190
rect 430 176 432 190
rect 458 176 460 190
rect 474 176 476 190
rect 531 176 533 190
rect 568 187 571 189
rect 575 187 582 189
rect 554 179 557 181
rect 561 179 568 181
rect 608 176 610 190
rect 639 176 641 190
rect 399 168 401 172
rect 430 168 432 172
rect 458 168 460 172
rect 474 168 476 172
rect 531 168 533 172
rect 608 168 610 172
rect 639 168 641 172
rect 376 145 383 147
rect 389 145 392 147
rect 395 145 398 147
rect 404 145 411 147
rect 416 145 423 147
rect 429 145 432 147
rect 435 145 438 147
rect 444 145 451 147
rect 557 144 559 151
rect 565 151 567 159
rect 565 145 567 147
rect 573 144 575 151
rect 585 145 592 147
rect 598 145 601 147
rect 604 145 607 147
rect 613 145 620 147
rect 625 145 632 147
rect 638 145 641 147
rect 644 145 647 147
rect 653 145 660 147
rect 512 137 519 139
rect 525 137 528 139
rect 531 137 534 139
rect 540 137 547 139
rect 557 137 559 140
rect 573 137 575 140
rect 472 132 474 135
rect 420 121 423 123
rect 426 121 440 123
rect 444 121 447 123
rect 585 123 592 125
rect 598 123 601 125
rect 604 123 607 125
rect 613 123 620 125
rect 625 123 632 125
rect 638 123 641 125
rect 644 123 647 125
rect 653 123 660 125
rect 472 107 474 121
rect 497 114 499 121
rect 497 105 499 108
rect 472 99 474 103
rect 497 99 499 102
rect 381 95 385 97
rect 389 95 403 97
rect 414 95 417 97
rect 591 96 595 98
rect 599 96 613 98
rect 624 96 627 98
rect 497 86 499 93
rect 550 92 552 95
rect 566 92 568 95
rect 550 67 552 81
rect 566 67 568 81
rect 630 66 634 68
rect 638 66 652 68
rect 663 66 666 68
rect 550 59 552 63
rect 566 59 568 63
<< polycontact >>
rect 473 380 477 384
rect 380 362 384 366
rect 411 362 415 366
rect 459 372 463 376
rect 503 372 507 376
rect 571 380 575 384
rect 445 364 449 368
rect 483 358 487 362
rect 503 356 507 360
rect 585 372 589 376
rect 540 362 544 366
rect 561 364 565 368
rect 630 362 634 366
rect 599 358 603 362
rect 661 362 665 366
rect 459 350 463 354
rect 561 348 565 352
rect 585 350 589 354
rect 473 342 477 346
rect 361 330 365 334
rect 392 330 396 334
rect 401 330 405 334
rect 432 330 436 334
rect 611 330 615 334
rect 642 330 646 334
rect 651 330 655 334
rect 682 330 686 334
rect 473 314 477 318
rect 361 308 365 312
rect 392 308 396 312
rect 401 308 405 312
rect 432 308 436 312
rect 487 322 491 326
rect 495 314 499 318
rect 519 316 523 320
rect 550 316 554 320
rect 571 315 575 319
rect 585 323 589 327
rect 593 315 597 319
rect 611 308 615 312
rect 642 308 646 312
rect 651 308 655 312
rect 682 308 686 312
rect 378 281 382 285
rect 465 284 469 288
rect 487 284 491 288
rect 503 284 507 288
rect 563 285 567 289
rect 585 285 589 289
rect 601 285 605 289
rect 628 281 632 285
rect 473 261 477 265
rect 495 261 499 265
rect 417 251 421 255
rect 667 251 671 255
rect 565 240 569 244
rect 581 240 585 244
rect 554 197 558 201
rect 395 179 399 183
rect 426 179 430 183
rect 460 179 464 183
rect 476 179 480 183
rect 533 179 537 183
rect 578 183 582 187
rect 604 179 608 183
rect 564 175 568 179
rect 635 179 639 183
rect 376 147 380 151
rect 407 147 411 151
rect 416 147 420 151
rect 447 147 451 151
rect 553 147 557 151
rect 567 155 571 159
rect 575 147 579 151
rect 585 147 589 151
rect 616 147 620 151
rect 625 147 629 151
rect 656 147 660 151
rect 512 133 516 137
rect 543 133 547 137
rect 429 123 433 127
rect 585 125 589 129
rect 616 125 620 129
rect 625 125 629 129
rect 656 125 660 129
rect 468 110 472 114
rect 499 117 503 121
rect 392 97 396 101
rect 602 98 606 102
rect 499 86 503 90
rect 546 70 550 74
rect 562 70 566 74
rect 641 68 645 72
<< polynplus >>
rect 384 355 386 356
rect 415 355 417 356
rect 538 355 540 356
rect 634 355 636 356
rect 665 355 667 356
rect 485 314 487 315
rect 583 315 585 316
rect 477 310 479 311
rect 493 310 495 311
rect 575 311 577 312
rect 591 311 593 312
rect 371 279 372 281
rect 621 279 622 281
rect 477 268 479 269
rect 493 268 495 269
rect 410 249 411 251
rect 660 249 661 251
rect 569 233 571 234
rect 585 233 587 234
rect 399 172 401 173
rect 430 172 432 173
rect 458 172 460 173
rect 474 172 476 173
rect 531 172 533 173
rect 608 172 610 173
rect 639 172 641 173
rect 565 147 567 148
rect 557 143 559 144
rect 573 143 575 144
rect 472 103 474 104
rect 385 95 386 97
rect 595 96 596 98
rect 550 63 552 64
rect 566 63 568 64
rect 634 66 635 68
<< metal1 >>
rect 371 395 429 396
rect 371 391 383 395
rect 387 391 414 395
rect 418 391 429 395
rect 371 390 429 391
rect 379 384 383 390
rect 410 384 414 390
rect 402 362 411 366
rect 379 351 383 355
rect 378 350 384 351
rect 378 346 379 350
rect 383 346 384 350
rect 378 345 384 346
rect 402 342 406 362
rect 410 351 414 355
rect 409 350 415 351
rect 409 346 410 350
rect 414 346 415 350
rect 409 345 415 346
rect 435 347 439 442
rect 444 395 511 396
rect 444 391 472 395
rect 476 391 511 395
rect 444 390 511 391
rect 527 390 552 396
rect 558 390 604 396
rect 621 395 679 396
rect 621 391 633 395
rect 637 391 664 395
rect 668 391 679 395
rect 621 390 679 391
rect 452 369 456 390
rect 466 377 470 390
rect 480 385 484 390
rect 541 384 545 390
rect 484 373 496 377
rect 564 385 568 390
rect 578 377 582 390
rect 480 365 496 369
rect 533 366 537 373
rect 568 369 572 377
rect 592 369 596 390
rect 629 384 633 390
rect 660 384 664 390
rect 466 361 470 365
rect 496 361 500 365
rect 526 362 537 366
rect 544 362 554 366
rect 435 343 445 347
rect 333 338 406 342
rect 353 320 357 338
rect 392 334 405 338
rect 441 334 445 343
rect 452 334 456 357
rect 476 349 480 357
rect 466 334 470 349
rect 480 334 484 341
rect 496 334 500 349
rect 441 330 500 334
rect 353 316 405 320
rect 480 319 484 330
rect 526 327 530 362
rect 533 359 537 362
rect 541 349 545 355
rect 540 348 546 349
rect 540 344 541 348
rect 545 344 546 348
rect 540 343 546 344
rect 550 331 554 362
rect 578 361 582 365
rect 652 362 661 366
rect 682 362 729 366
rect 568 353 572 357
rect 568 331 572 341
rect 578 334 582 349
rect 592 334 596 357
rect 629 351 633 355
rect 628 350 634 351
rect 628 346 629 350
rect 633 346 634 350
rect 628 345 634 346
rect 652 342 656 362
rect 660 351 664 355
rect 659 350 665 351
rect 659 346 660 350
rect 664 346 665 350
rect 659 345 665 346
rect 682 342 686 362
rect 652 340 694 342
rect 651 338 694 340
rect 578 331 596 334
rect 543 330 596 331
rect 642 334 655 338
rect 543 327 582 330
rect 578 320 582 327
rect 690 320 694 338
rect 361 312 365 316
rect 401 312 405 316
rect 488 311 492 315
rect 484 307 488 311
rect 374 301 383 305
rect 414 301 423 305
rect 472 303 476 307
rect 496 303 500 307
rect 360 285 371 286
rect 360 281 361 285
rect 365 282 371 285
rect 378 285 382 301
rect 406 286 412 294
rect 365 281 366 282
rect 400 282 412 286
rect 360 280 366 281
rect 406 278 407 282
rect 411 278 412 282
rect 406 267 412 278
rect 398 256 404 257
rect 398 252 399 256
rect 403 252 410 256
rect 417 255 421 301
rect 472 299 500 303
rect 472 295 476 299
rect 488 295 492 299
rect 458 291 464 295
rect 496 295 500 299
rect 445 256 451 264
rect 458 260 462 291
rect 480 280 484 291
rect 472 276 500 280
rect 472 272 476 276
rect 480 275 484 276
rect 496 272 500 276
rect 484 261 488 272
rect 398 251 404 252
rect 439 252 451 256
rect 445 248 446 252
rect 450 248 451 252
rect 414 244 428 248
rect 417 233 421 244
rect 445 237 451 248
rect 519 233 523 316
rect 532 315 541 319
rect 534 244 538 315
rect 586 312 590 316
rect 611 316 694 320
rect 611 312 615 316
rect 582 308 586 312
rect 651 312 655 316
rect 570 304 574 308
rect 594 304 598 308
rect 570 300 606 304
rect 624 301 633 305
rect 664 301 673 305
rect 570 296 574 300
rect 586 296 590 300
rect 602 296 606 300
rect 556 292 562 296
rect 556 281 560 292
rect 578 281 582 292
rect 594 281 598 292
rect 610 285 621 286
rect 556 277 598 281
rect 610 281 611 285
rect 615 282 621 285
rect 628 285 632 301
rect 656 286 662 294
rect 615 281 616 282
rect 650 282 662 286
rect 610 280 616 281
rect 656 278 657 282
rect 661 278 662 282
rect 556 273 599 274
rect 556 269 568 273
rect 572 269 584 273
rect 588 269 599 273
rect 556 268 599 269
rect 564 262 568 268
rect 580 262 584 268
rect 656 267 662 278
rect 648 256 654 257
rect 648 252 649 256
rect 653 252 660 256
rect 667 255 671 301
rect 695 256 701 264
rect 648 251 654 252
rect 689 252 701 256
rect 572 244 576 251
rect 588 244 592 251
rect 695 248 696 252
rect 700 248 701 252
rect 534 240 565 244
rect 572 240 581 244
rect 588 240 603 244
rect 572 237 576 240
rect 588 237 592 240
rect 417 229 523 233
rect 564 227 568 233
rect 580 227 584 233
rect 563 226 569 227
rect 563 222 564 226
rect 568 222 569 226
rect 563 221 569 222
rect 579 226 585 227
rect 579 222 580 226
rect 584 222 585 226
rect 579 221 585 222
rect 599 225 603 240
rect 695 237 701 248
rect 599 221 688 225
rect 386 212 488 213
rect 386 208 398 212
rect 402 208 429 212
rect 433 208 457 212
rect 461 208 473 212
rect 477 208 488 212
rect 386 207 488 208
rect 520 212 545 213
rect 520 208 530 212
rect 534 208 545 212
rect 520 207 545 208
rect 551 212 583 213
rect 551 208 564 212
rect 568 208 583 212
rect 551 207 583 208
rect 595 212 653 213
rect 595 208 607 212
rect 611 208 638 212
rect 642 208 653 212
rect 595 207 653 208
rect 394 201 398 207
rect 425 201 429 207
rect 461 201 465 207
rect 477 201 481 207
rect 534 201 538 207
rect 561 202 565 207
rect 571 194 575 207
rect 603 201 607 207
rect 634 201 638 207
rect 469 183 473 190
rect 526 183 530 190
rect 561 189 565 190
rect 557 186 565 189
rect 416 179 426 183
rect 464 179 473 183
rect 480 179 495 183
rect 394 167 398 172
rect 393 166 399 167
rect 393 162 394 166
rect 398 162 399 166
rect 393 161 399 162
rect 416 158 420 179
rect 469 176 473 179
rect 425 166 429 172
rect 461 166 465 172
rect 477 166 481 172
rect 424 165 430 166
rect 424 161 425 165
rect 429 161 430 165
rect 424 160 430 161
rect 460 165 466 166
rect 460 161 461 165
rect 465 161 466 165
rect 460 160 466 161
rect 476 165 482 166
rect 476 161 477 165
rect 481 161 482 165
rect 476 160 482 161
rect 333 155 420 158
rect 407 151 420 155
rect 389 140 398 144
rect 459 143 486 144
rect 373 102 379 103
rect 373 98 374 102
rect 378 98 385 102
rect 392 101 396 140
rect 459 139 471 143
rect 475 139 486 143
rect 459 138 486 139
rect 410 128 416 129
rect 449 128 455 134
rect 410 124 411 128
rect 415 124 422 128
rect 410 123 416 124
rect 444 124 455 128
rect 449 120 450 124
rect 454 120 455 124
rect 467 132 471 138
rect 491 129 495 179
rect 519 179 530 183
rect 537 179 547 183
rect 519 144 523 179
rect 526 176 530 179
rect 534 166 538 172
rect 533 165 539 166
rect 533 161 534 165
rect 538 161 539 165
rect 533 160 539 161
rect 543 165 547 179
rect 557 172 561 174
rect 571 172 575 182
rect 626 179 635 183
rect 664 179 711 183
rect 557 168 575 172
rect 603 168 607 172
rect 566 165 570 168
rect 543 162 570 165
rect 602 167 608 168
rect 602 163 603 167
rect 607 163 608 167
rect 602 162 608 163
rect 543 161 564 162
rect 543 148 547 161
rect 560 152 564 161
rect 626 159 630 179
rect 634 168 638 172
rect 633 167 639 168
rect 633 163 634 167
rect 638 163 639 167
rect 633 162 639 163
rect 664 159 668 179
rect 626 157 668 159
rect 625 155 668 157
rect 536 144 547 148
rect 568 144 572 148
rect 616 151 629 155
rect 564 140 568 144
rect 525 132 534 136
rect 552 136 556 140
rect 576 136 580 140
rect 664 137 668 155
rect 552 135 580 136
rect 491 125 511 129
rect 426 116 440 120
rect 420 102 426 110
rect 429 106 433 116
rect 449 110 455 120
rect 475 114 479 121
rect 459 110 468 114
rect 475 110 492 114
rect 459 106 463 110
rect 475 107 479 110
rect 429 102 463 106
rect 373 97 379 98
rect 414 98 426 102
rect 420 94 421 98
rect 425 94 426 98
rect 389 90 403 94
rect 392 28 396 90
rect 420 83 426 94
rect 459 87 463 102
rect 500 106 504 108
rect 507 106 511 125
rect 467 97 471 103
rect 500 102 511 106
rect 500 99 504 102
rect 466 96 472 97
rect 466 92 467 96
rect 471 92 472 96
rect 466 91 472 92
rect 483 93 492 97
rect 483 87 487 93
rect 459 83 487 87
rect 527 74 531 132
rect 552 131 564 135
rect 568 131 580 135
rect 552 130 580 131
rect 585 133 668 137
rect 585 129 589 133
rect 625 129 629 133
rect 598 118 607 122
rect 638 118 647 122
rect 537 103 580 104
rect 537 99 549 103
rect 553 99 565 103
rect 569 99 580 103
rect 537 98 580 99
rect 583 103 589 104
rect 583 99 584 103
rect 588 99 595 103
rect 602 102 606 118
rect 630 103 636 111
rect 583 98 589 99
rect 624 99 636 103
rect 545 92 549 98
rect 561 92 565 98
rect 630 95 631 99
rect 635 95 636 99
rect 630 84 636 95
rect 553 74 557 81
rect 569 74 573 81
rect 527 70 546 74
rect 553 70 562 74
rect 569 70 580 74
rect 553 67 557 70
rect 569 67 573 70
rect 455 28 459 64
rect 545 57 549 63
rect 561 57 565 63
rect 544 56 550 57
rect 544 52 545 56
rect 549 52 550 56
rect 544 51 550 52
rect 560 56 566 57
rect 560 52 561 56
rect 565 52 566 56
rect 560 51 566 52
rect 576 28 580 70
rect 622 73 628 74
rect 622 69 623 73
rect 627 69 634 73
rect 641 72 645 118
rect 669 73 675 81
rect 622 68 628 69
rect 663 69 675 73
rect 669 65 670 69
rect 674 65 675 69
rect 669 54 675 65
rect 689 28 693 128
<< m2contact >>
rect 688 220 694 226
rect 688 128 694 134
rect 454 64 460 70
<< metal2 >>
rect 387 366 391 373
rect 637 366 641 373
rect 387 362 399 366
rect 387 359 391 362
rect 395 342 399 362
rect 637 362 649 366
rect 637 359 641 362
rect 645 342 649 362
rect 353 338 429 342
rect 353 316 357 338
rect 385 335 389 338
rect 425 335 429 338
rect 635 338 694 342
rect 635 335 639 338
rect 675 335 679 338
rect 690 320 694 338
rect 370 316 429 320
rect 620 316 694 320
rect 370 313 374 316
rect 425 313 429 316
rect 375 274 389 278
rect 377 233 381 274
rect 550 233 554 316
rect 620 313 624 316
rect 675 313 679 316
rect 664 244 678 248
rect 377 229 554 233
rect 667 218 671 244
rect 507 214 671 218
rect 402 183 406 190
rect 453 183 457 190
rect 402 179 413 183
rect 402 176 406 179
rect 410 159 413 179
rect 445 179 457 183
rect 445 160 449 179
rect 453 176 457 179
rect 383 156 429 159
rect 445 156 459 160
rect 383 152 387 156
rect 393 155 419 156
rect 425 152 429 156
rect 455 70 459 156
rect 507 137 511 214
rect 611 183 615 190
rect 611 179 623 183
rect 611 176 615 179
rect 619 159 623 179
rect 609 156 668 159
rect 609 155 643 156
rect 649 155 668 156
rect 609 152 613 155
rect 649 152 653 155
rect 664 137 668 155
rect 507 133 512 137
rect 594 134 668 137
rect 689 134 693 220
rect 594 133 643 134
rect 649 133 668 134
rect 594 130 598 133
rect 649 130 653 133
rect 599 91 613 95
rect 503 86 519 90
rect 515 49 519 86
rect 602 49 606 91
rect 515 45 606 49
<< metal3 >>
rect 514 389 609 393
rect 438 380 473 384
rect 438 376 442 380
rect 438 372 459 376
rect 333 362 380 366
rect 370 342 374 362
rect 353 338 374 342
rect 353 319 357 338
rect 438 327 442 372
rect 459 340 463 350
rect 514 340 518 389
rect 605 362 609 389
rect 603 358 609 362
rect 459 336 518 340
rect 414 323 423 327
rect 429 323 477 327
rect 353 318 405 319
rect 353 315 414 318
rect 385 313 389 315
rect 410 313 414 315
rect 454 288 458 323
rect 473 318 477 323
rect 499 314 503 336
rect 585 335 589 350
rect 559 331 589 335
rect 559 319 563 331
rect 605 327 609 358
rect 620 362 630 366
rect 620 342 624 362
rect 620 338 729 342
rect 589 323 618 327
rect 624 323 633 327
rect 690 319 694 338
rect 559 315 571 319
rect 635 316 694 319
rect 559 304 563 315
rect 635 313 639 316
rect 660 313 664 316
rect 548 300 563 304
rect 454 284 465 288
rect 512 233 516 238
rect 548 233 552 300
rect 512 229 552 233
rect 548 218 552 229
rect 548 214 590 218
rect 333 179 395 183
rect 578 179 582 183
rect 586 179 590 214
rect 386 159 390 179
rect 578 175 590 179
rect 594 179 604 183
rect 578 161 582 175
rect 572 159 584 161
rect 386 155 402 159
rect 571 157 584 159
rect 571 155 575 157
rect 398 152 402 155
rect 581 144 584 157
rect 594 159 598 179
rect 594 155 711 159
rect 581 140 592 144
rect 598 140 607 144
rect 625 136 637 137
rect 664 136 668 155
rect 609 134 668 136
rect 609 133 628 134
rect 634 133 668 134
rect 609 130 613 133
rect 634 130 638 133
<< metal4 >>
rect 514 389 609 393
rect 514 376 518 389
rect 605 384 609 389
rect 575 380 609 384
rect 605 376 609 380
rect 507 372 518 376
rect 589 372 609 376
rect 438 364 445 368
rect 555 364 561 368
rect 438 332 442 364
rect 438 328 491 332
rect 505 330 516 334
rect 374 323 383 327
rect 376 319 379 323
rect 438 319 442 328
rect 487 326 491 328
rect 359 316 442 319
rect 512 289 516 330
rect 555 304 559 364
rect 605 320 609 372
rect 664 324 673 327
rect 667 323 673 324
rect 667 320 671 323
rect 605 319 671 320
rect 597 316 671 319
rect 597 315 609 316
rect 548 300 559 304
rect 605 304 609 315
rect 605 300 615 304
rect 548 289 552 300
rect 611 289 615 300
rect 512 288 519 289
rect 507 285 519 288
rect 523 285 563 289
rect 605 286 615 289
rect 507 284 516 285
rect 512 265 516 284
rect 499 261 516 265
rect 548 218 552 285
rect 625 274 639 278
rect 628 218 632 274
rect 507 214 632 218
rect 507 129 511 214
rect 586 179 590 214
rect 568 175 590 179
rect 580 151 583 175
rect 579 147 584 151
rect 581 136 584 147
rect 638 140 647 144
rect 641 136 645 140
rect 581 133 645 136
rect 543 129 547 133
rect 507 125 547 129
<< m345contact >>
rect 511 238 517 244
<< m5contact >>
rect 499 329 505 335
<< metal5 >>
rect 418 366 422 373
rect 668 366 672 373
rect 418 362 436 366
rect 668 362 686 366
rect 418 359 422 362
rect 432 342 436 362
rect 487 358 492 362
rect 353 338 436 342
rect 353 320 357 338
rect 361 334 365 338
rect 432 334 436 338
rect 473 329 477 342
rect 488 334 492 358
rect 507 356 516 360
rect 668 359 672 362
rect 488 330 499 334
rect 454 325 477 329
rect 353 316 436 320
rect 392 312 396 316
rect 432 312 436 316
rect 454 265 458 325
rect 487 282 491 284
rect 512 282 516 356
rect 555 348 561 352
rect 555 304 559 348
rect 682 342 686 362
rect 611 338 694 342
rect 611 334 615 338
rect 682 334 686 338
rect 690 320 694 338
rect 642 316 694 320
rect 642 312 646 316
rect 690 312 694 316
rect 686 308 694 312
rect 487 278 516 282
rect 454 261 473 265
rect 454 222 458 261
rect 512 244 516 278
rect 546 300 559 304
rect 546 282 550 300
rect 585 282 589 285
rect 546 278 589 282
rect 454 218 497 222
rect 433 183 437 190
rect 433 179 451 183
rect 433 176 437 179
rect 447 159 451 179
rect 376 155 451 159
rect 493 157 497 218
rect 546 201 550 278
rect 546 197 554 201
rect 546 157 550 197
rect 642 183 646 190
rect 642 179 660 183
rect 642 176 646 179
rect 656 159 660 179
rect 376 151 380 155
rect 447 151 451 155
rect 461 153 557 157
rect 429 140 438 144
rect 430 136 434 140
rect 461 136 465 153
rect 553 151 557 153
rect 585 155 668 159
rect 585 151 589 155
rect 656 151 660 155
rect 664 136 668 155
rect 429 132 465 136
rect 616 133 668 136
rect 429 127 433 132
rect 616 129 620 133
rect 664 129 668 133
rect 660 125 668 129
rect 503 117 519 121
rect 515 49 519 117
rect 638 61 652 65
rect 641 49 645 61
rect 515 45 645 49
<< labels >>
rlabel pdcontact 380 377 382 379 1 vdd
rlabel nwell 534 385 536 387 1 vdd
rlabel ndcontact 505 292 507 294 1 gnd
rlabel nwell 403 375 405 377 1 vdd
rlabel pdcontact 411 377 413 379 1 vdd
rlabel ndcontact 465 292 467 294 1 gnd
rlabel ndcontact 481 269 483 271 1 gnd
rlabel ndcontact 489 269 491 271 1 gnd
rlabel ndcontact 497 269 499 271 1 node14
rlabel ndcontact 473 269 475 271 1 node14
rlabel ndcontact 481 292 483 294 1 node14
rlabel ndcontact 497 292 499 294 1 node13
rlabel ndcontact 489 292 491 294 1 node13
rlabel ndcontact 473 292 475 294 1 node13
rlabel ndcontact 473 308 475 310 1 node13
rlabel ndcontact 497 308 499 310 1 node13
rlabel ndcontact 489 308 491 310 1 node12
rlabel ndcontact 481 308 483 310 1 node12
rlabel ndcontact 489 316 491 318 1 node12
rlabel pdcontact 481 342 483 344 1 C4
rlabel pdcontact 481 350 483 352 1 node11
rlabel pdcontact 477 358 479 360 1 node11
rlabel pdcontact 497 358 499 360 1 node10
rlabel pdcontact 477 366 479 368 1 node10
rlabel pdcontact 497 366 499 368 1 node10
rlabel pdcontact 497 374 499 376 1 node9
rlabel pdcontact 481 374 483 376 1 node9
rlabel pdcontact 467 358 469 360 1 node8
rlabel pdcontact 467 366 469 368 1 node8
rlabel nwell 493 381 495 383 1 vdd
rlabel pdcontact 481 382 483 384 1 vdd
rlabel pdcontact 467 374 469 376 1 vdd
rlabel pdcontact 453 366 455 368 1 vdd
rlabel polycontact 551 317 553 319 1 P_not4
rlabel polycontact 520 317 522 319 1 P4
rlabel pdcontact 433 253 435 255 1 vdd
rlabel ndcontact 411 245 413 247 1 P4
rlabel pdcontact 432 245 434 247 1 P4
rlabel pdcontact 393 275 395 277 1 P_not4
rlabel ndcontact 372 275 374 277 1 P_not4
rlabel pdcontact 393 283 395 285 1 vdd
rlabel polycontact 379 282 381 284 1 P_4
rlabel ndcontact 385 302 387 304 1 P_4
rlabel ndcontact 370 302 372 304 1 P_4
rlabel polycontact 418 252 420 254 1 P_not_4
rlabel ndcontact 425 302 427 304 1 P_not_4
rlabel ndcontact 410 302 412 304 1 P_not_4
rlabel polycontact 488 285 490 287 1 G_2
rlabel polycontact 466 285 468 287 1 K_4
rlabel polycontact 496 262 498 264 1 K_2
rlabel polycontact 474 262 476 264 1 G_1
rlabel polycontact 474 315 476 317 1 K_4
rlabel polycontact 496 315 498 317 1 G_3
rlabel ndcontact 481 316 483 318 1 C4
rlabel pdcontact 453 358 455 360 1 C4
rlabel pdcontact 467 350 469 352 1 C4
rlabel pdcontact 497 350 499 352 1 C4
rlabel polycontact 474 343 476 345 1 G_1
rlabel polycontact 504 357 506 359 1 G_2
rlabel polycontact 484 359 486 361 1 K_2
rlabel polycontact 504 373 506 375 1 K_3
rlabel ndcontact 370 332 372 334 1 vdd
rlabel polycontact 381 363 383 365 1 B4
rlabel ndcontact 385 310 387 312 1 B4
rlabel ndcontact 410 310 412 312 1 B4
rlabel pdcontact 388 377 390 379 1 B_not4
rlabel ndcontact 388 356 390 358 1 B_not4
rlabel ndcontact 385 332 387 334 1 B_not4
rlabel ndcontact 425 332 427 334 1 B_not4
rlabel ndcontact 425 310 427 312 1 B_not4
rlabel ndcontact 370 310 372 312 1 B_not4
rlabel polycontact 412 363 414 365 1 A4
rlabel polycontact 402 331 404 333 1 A4
rlabel polycontact 393 331 395 333 1 A4
rlabel polycontact 402 309 404 311 1 A4
rlabel polycontact 362 309 364 311 1 A4
rlabel pdcontact 419 378 421 380 1 A_not4
rlabel ndcontact 419 356 421 358 1 A_not4
rlabel polycontact 433 331 435 333 1 A_not4
rlabel polycontact 362 331 364 333 1 A_not4
rlabel polycontact 393 309 395 311 1 A_not4
rlabel polycontact 433 309 435 311 1 A_not4
rlabel ndcontact 410 332 412 334 1 gnd
rlabel ndcontact 411 356 413 358 1 gnd
rlabel ndcontact 380 356 382 358 1 gnd
rlabel ndcontact 372 283 374 285 1 gnd
rlabel ndcontact 411 253 413 255 1 gnd
rlabel ndcontact 370 324 372 326 1 G_4
rlabel ndcontact 385 324 387 326 1 G_4
rlabel ndcontact 410 324 412 326 1 K_4
rlabel ndcontact 425 324 427 326 1 K_4
rlabel polycontact 446 365 448 367 5 G_4
rlabel polycontact 488 323 490 325 1 G_4
rlabel polycontact 460 351 462 353 1 G_3
rlabel polycontact 474 381 476 383 1 K_4
rlabel polycontact 460 373 462 375 1 K_4
rlabel nwell 584 365 586 367 1 vdd
rlabel pdcontact 581 255 583 257 1 vdd
rlabel pdcontact 589 256 591 258 1 S4
rlabel ndcontact 589 234 591 236 1 S4
rlabel polycontact 582 241 584 243 1 S_4
rlabel pdcontact 573 256 575 258 1 S_4
rlabel ndcontact 573 234 575 236 1 S_4
rlabel polycontact 566 241 568 243 1 sum4
rlabel ndcontact 543 316 545 318 1 sum4
rlabel ndcontact 528 316 530 318 1 sum4
rlabel pdcontact 534 377 536 379 1 C_not3
rlabel ndcontact 534 356 536 358 1 C_not3
rlabel ndcontact 528 324 530 326 1 C_not3
rlabel polycontact 541 363 543 365 1 C3
rlabel ndcontact 543 324 545 326 1 C3
rlabel ndcontact 603 293 605 295 1 node7
rlabel ndcontact 587 293 589 295 1 node7
rlabel ndcontact 571 293 573 295 1 node7
rlabel ndcontact 595 309 597 311 1 node7
rlabel ndcontact 571 309 573 311 1 node7
rlabel ndcontact 579 309 581 311 1 node6
rlabel ndcontact 587 309 589 311 1 node6
rlabel ndcontact 587 317 589 319 1 node6
rlabel ndcontact 579 317 581 319 1 C3
rlabel pdcontact 593 358 595 360 1 C3
rlabel pdcontact 569 342 571 344 1 C3
rlabel pdcontact 579 350 581 352 1 C3
rlabel pdcontact 579 358 581 360 1 node5
rlabel pdcontact 579 366 581 368 1 node5
rlabel pdcontact 569 350 571 352 1 node4
rlabel pdcontact 569 358 571 360 1 node4
rlabel pdcontact 569 366 571 368 1 node3
rlabel pdcontact 565 374 567 376 1 node3
rlabel polycontact 586 286 588 288 1 G_1
rlabel polycontact 564 286 566 288 1 K_2
rlabel polycontact 572 316 574 318 1 G_2
rlabel polycontact 586 324 588 326 1 G_3
rlabel polycontact 594 316 596 318 1 K_3
rlabel polycontact 600 359 602 361 1 G_3
rlabel polycontact 562 365 564 367 1 K_2
rlabel polycontact 562 349 564 351 1 G_1
rlabel polycontact 586 351 588 353 1 G_2
rlabel ndcontact 542 356 544 358 1 gnd
rlabel ndcontact 595 293 597 295 1 gnd
rlabel ndcontact 579 293 581 295 1 gnd
rlabel ndcontact 563 293 565 295 1 gnd
rlabel ndcontact 581 234 583 236 1 gnd
rlabel ndcontact 565 234 567 236 1 gnd
rlabel ndcontact 630 356 632 358 1 gnd
rlabel ndcontact 661 356 663 358 1 gnd
rlabel ndcontact 661 253 663 255 1 gnd
rlabel ndcontact 622 283 624 285 1 gnd
rlabel polycontact 668 252 670 254 1 P_not_3
rlabel polycontact 629 282 631 284 1 P_3
rlabel ndcontact 675 302 677 304 1 P_not_3
rlabel ndcontact 660 302 662 304 1 P_not_3
rlabel ndcontact 635 302 637 304 1 P_3
rlabel ndcontact 620 302 622 304 1 P_3
rlabel polycontact 586 373 588 375 1 K_3
rlabel polycontact 572 381 574 383 1 K_3
rlabel polycontact 602 286 604 288 1 K_3
rlabel ndcontact 675 324 677 326 1 K_3
rlabel ndcontact 660 324 662 326 1 K_3
rlabel ndcontact 635 324 637 326 1 G_3
rlabel ndcontact 620 324 622 326 1 G_3
rlabel polycontact 683 309 685 311 1 A_not3
rlabel polycontact 643 309 645 311 1 A_not3
rlabel polycontact 612 331 614 333 1 A_not3
rlabel polycontact 683 331 685 333 1 A_not3
rlabel ndcontact 669 356 671 358 1 A_not3
rlabel pdcontact 669 377 671 379 1 A_not3
rlabel ndcontact 660 332 662 334 1 gnd
rlabel polycontact 612 309 614 311 1 A3
rlabel polycontact 652 309 654 311 1 A3
rlabel polycontact 643 331 645 333 1 A3
rlabel polycontact 652 331 654 333 1 A3
rlabel polycontact 662 363 664 365 1 A3
rlabel ndcontact 620 310 622 312 1 B_not3
rlabel ndcontact 675 310 677 312 1 B_not3
rlabel ndcontact 675 332 677 334 1 B_not3
rlabel ndcontact 635 332 637 334 1 B_not3
rlabel ndcontact 638 356 640 358 1 B_not3
rlabel pdcontact 638 377 640 379 1 B_not3
rlabel pdcontact 565 255 567 257 1 vdd
rlabel pdcontact 542 377 544 379 1 vdd
rlabel pdcontact 565 382 567 384 1 vdd
rlabel pdcontact 579 374 581 376 1 vdd
rlabel pdcontact 593 366 595 368 1 vdd
rlabel pdcontact 682 253 684 255 1 vdd
rlabel pdcontact 643 283 645 285 1 vdd
rlabel pdcontact 661 377 663 379 1 vdd
rlabel pdcontact 630 377 632 379 1 vdd
rlabel ndcontact 635 310 637 312 1 B3
rlabel ndcontact 660 310 662 312 1 B3
rlabel polycontact 631 363 633 365 1 B3
rlabel pdcontact 643 275 645 277 1 P_not3
rlabel ndcontact 622 275 624 277 1 P_not3
rlabel pdcontact 682 245 684 247 1 P3
rlabel ndcontact 661 245 663 247 1 P3
rlabel ndcontact 620 332 622 334 1 vdd
rlabel polycontact 504 285 506 287 1 K_2
rlabel polycontact 500 118 502 120 1 P2
rlabel ndcontact 476 104 478 106 1 C_not1
rlabel pdcontact 476 125 478 128 1 C_not1
rlabel polycontact 544 134 546 136 1 P_not3
rlabel polycontact 513 134 515 136 1 P3
rlabel ndcontact 634 149 636 151 1 gnd
rlabel ndcontact 635 173 637 175 1 gnd
rlabel pdcontact 570 85 572 87 1 S3
rlabel ndcontact 570 64 572 66 1 S3
rlabel ndcontact 554 64 556 66 1 s_3
rlabel pdcontact 554 85 556 87 1 s_3
rlabel polycontact 563 71 565 73 1 s_3
rlabel polycontact 547 71 549 73 1 sum3
rlabel ndcontact 536 133 538 135 1 sum3
rlabel ndcontact 521 133 523 135 1 sum3
rlabel ndcontact 535 173 537 175 1 gnd
rlabel pdcontact 535 194 537 196 1 vdd
rlabel pdcontact 527 194 529 196 1 C_not2
rlabel ndcontact 527 173 529 175 1 C_not2
rlabel ndcontact 521 141 523 143 1 C_not2
rlabel ndcontact 536 141 538 143 1 C2
rlabel polycontact 534 180 536 182 1 C2
rlabel ndcontact 553 141 555 143 1 gnd
rlabel ndcontact 577 141 579 143 1 gnd
rlabel ndcontact 561 141 563 143 1 node1
rlabel ndcontact 569 141 571 143 1 node1
rlabel ndcontact 569 149 571 151 1 node1
rlabel ndcontact 561 149 563 151 1 C2
rlabel pdcontact 572 183 574 185 1 C2
rlabel pdcontact 558 175 560 177 1 C2
rlabel pdcontact 572 191 574 193 1 vdd
rlabel pdcontact 562 199 564 201 1 vdd
rlabel pdcontact 558 183 560 185 1 node2
rlabel pdcontact 562 191 564 193 1 node2
rlabel ndcontact 562 64 564 66 1 gnd
rlabel ndcontact 546 64 548 66 1 gnd
rlabel ndcontact 596 100 598 102 1 gnd
rlabel ndcontact 635 70 637 72 1 gnd
rlabel pdcontact 617 92 619 94 1 P_not2
rlabel ndcontact 596 92 598 94 1 P_not2
rlabel polycontact 603 99 605 101 1 P_2
rlabel pdcontact 656 62 658 64 1 P2
rlabel ndcontact 635 62 637 64 1 P2
rlabel polycontact 642 69 644 71 1 P_not_2
rlabel ndcontact 649 119 651 121 1 P_not_2
rlabel ndcontact 634 119 636 121 1 P_not_2
rlabel ndcontact 609 119 611 121 1 P_2
rlabel ndcontact 594 119 596 121 1 P_2
rlabel polycontact 565 176 567 178 1 K_2
rlabel polycontact 576 148 578 150 1 K_2
rlabel ndcontact 649 141 651 143 1 K_2
rlabel ndcontact 634 141 636 143 1 K_2
rlabel polycontact 579 184 581 186 1 G_2
rlabel polycontact 568 156 570 158 1 G_2
rlabel ndcontact 609 141 611 143 1 G_2
rlabel ndcontact 594 141 596 143 1 G_2
rlabel ndcontact 594 149 596 151 1 vdd
rlabel polycontact 657 126 659 128 1 A_not2
rlabel polycontact 617 126 619 128 1 A_not2
rlabel polycontact 586 148 588 150 1 A_not2
rlabel polycontact 657 148 659 150 1 A_not2
rlabel ndcontact 643 173 645 175 1 A_not2
rlabel pdcontact 643 195 645 197 1 A_not2
rlabel polycontact 586 126 588 128 1 A2
rlabel polycontact 626 126 628 128 1 A2
rlabel polycontact 617 148 619 150 1 A2
rlabel polycontact 626 148 628 150 1 A2
rlabel polycontact 636 180 638 182 1 A2
rlabel ndcontact 594 127 596 129 1 B_not2
rlabel ndcontact 649 127 651 129 1 B_not2
rlabel ndcontact 649 149 651 151 1 B_not2
rlabel ndcontact 609 149 611 151 1 B_not2
rlabel metal2 612 180 614 182 1 B_not2
rlabel ndcontact 612 173 614 175 1 B_not2
rlabel pdcontact 612 194 614 196 1 B_not2
rlabel ndcontact 609 127 611 129 1 B2
rlabel ndcontact 634 127 636 129 1 B2
rlabel polycontact 605 180 607 182 1 B2
rlabel nwell 540 85 542 87 1 vdd
rlabel pdcontact 546 86 548 88 1 vdd
rlabel pdcontact 562 86 564 88 1 vdd
rlabel pdcontact 656 70 658 72 1 vdd
rlabel nwell 620 105 622 107 1 vdd
rlabel pdcontact 617 100 619 102 1 vdd
rlabel pdcontact 635 195 637 197 1 vdd
rlabel nwell 598 194 600 196 1 vdd
rlabel pdcontact 604 194 606 196 1 vdd
rlabel polycontact 554 148 556 150 1 G_1
rlabel polycontact 555 198 557 200 1 G_1
rlabel ndcontact 604 173 606 175 1 gnd
rlabel pdcontact 395 194 397 196 1 vdd
rlabel polycontact 396 180 398 182 1 B1
rlabel ndcontact 400 149 402 151 1 B1
rlabel pdcontact 403 195 405 197 1 B_not1
rlabel ndcontact 385 149 387 151 1 B_not1
rlabel ndcontact 425 149 427 151 1 B_not1
rlabel ndcontact 440 149 442 151 1 vdd
rlabel pdcontact 426 195 428 197 1 vdd
rlabel nwell 415 195 417 197 1 vdd
rlabel pdcontact 407 99 409 101 1 vdd
rlabel pdcontact 441 125 443 127 1 vdd
rlabel pdcontact 468 126 470 128 1 vdd
rlabel nwell 463 127 465 129 1 vdd
rlabel polycontact 427 180 429 182 1 A1
rlabel pdcontact 434 194 436 196 1 A_not1
rlabel ndcontact 434 173 436 175 1 A_not1
rlabel polycontact 377 148 379 150 1 A_not1
rlabel polycontact 448 148 450 150 1 A_not1
rlabel polycontact 408 148 410 150 1 A1
rlabel polycontact 417 148 419 150 1 A1
rlabel ndcontact 400 141 402 143 1 P_not1
rlabel ndcontact 385 141 387 143 1 P_not1
rlabel polycontact 393 98 395 100 1 P_not1
rlabel metal1 393 91 395 93 1 S1
rlabel ndcontact 386 91 388 93 1 S1
rlabel pdcontact 407 91 409 93 1 S1
rlabel ndcontact 425 141 427 143 1 G_1
rlabel ndcontact 440 141 442 143 1 G_1
rlabel polycontact 430 124 432 126 1 G_1
rlabel ndcontact 386 99 388 101 1 gnd
rlabel ndcontact 423 125 425 127 1 gnd
rlabel ndcontact 395 173 397 175 1 gnd
rlabel ndcontact 426 173 428 175 1 gnd
rlabel ndcontact 468 104 470 106 1 gnd
rlabel pdcontact 441 117 443 119 1 C1
rlabel ndcontact 423 117 425 119 1 C1
rlabel polycontact 469 111 471 113 1 C1
rlabel ndcontact 493 95 495 97 1 C1
rlabel ndcontact 493 110 495 112 1 C_not1
rlabel polycontact 500 87 502 89 1 P_not2
rlabel ndcontact 501 110 503 112 1 sum2
rlabel ndcontact 501 95 503 97 1 sum2
rlabel polycontact 477 180 479 182 1 sum2
rlabel ndcontact 478 173 480 175 1 gnd
rlabel ndcontact 462 173 464 175 1 gnd
rlabel ndcontact 470 173 472 175 1 S_2
rlabel pdcontact 470 194 472 196 1 S_2
rlabel polycontact 461 180 463 182 1 S_2
rlabel ndcontact 454 173 456 175 1 S2
rlabel pdcontact 454 195 456 197 1 S2
rlabel pdcontact 462 195 464 197 1 vdd
rlabel nwell 466 195 468 197 1 vdd
rlabel pdcontact 478 195 480 197 1 vdd
rlabel ndcontact 403 173 405 175 1 B_not1
<< end >>
